library IEEE;
use IEEE.STD_LOGIC_1164.all;
--use IEEE.std_logic_unsigned.all;
--use ieee.numeric_std.all;
--use ieee.std_logic_arith.all;



entity rec_object is
port 	(
		--////////////////////	Clock Input	 	////////////////////	
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		Record1Enable : in std_logic;
		--ObjectStartX	: in integer;
		--ObjectStartY 	: in integer;
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0) 
	);
end entity;

architecture behav of rec_object is 
constant StartX : integer := 285;   -- starting point
constant StartY : integer := 270;
constant object_X_size : integer := 60;
constant object_Y_size : integer := 60;
--constant R_high		: integer := 7;
--constant R_low		: integer := 5;
--constant G_high		: integer := 4;
--constant G_low		: integer := 2;
--constant B_high		: integer := 1;
--constant B_low		: integer := 0;


type object_form is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object : object_form := (
("000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000001111111100000000000000000000000000"),
("000000000000000000000111111111111111111000000000000000000000"),
("000000000000000000111111111111111111111111000000000000000000"),
("000000000000000011111111111111111111111111110000000000000000"),
("000000000000000111111111111111111111111111111000000000000000"),
("000000000000011111111111111111111111111111111110000000000000"),
("000000000000111111111111111111111111111111111111000000000000"),
("000000000001111111111111111111111111111111111111100000000000"),
("000000000011111111111111111111111111111111111111110000000000"),
("000000000111111111111111111111111111111111111111111000000000"),
("000000001111111111111111111111111111111111111111111100000000"),
("000000011111111111111111111111111111111111111111111110000000"),
("000000111111111111111111111111111111111111111111111111000000"),
("000000111111111111111111111111111111111111111111111111100000"),
("000001111111111111111111111111111111111111111111111111100000"),
("000011111111111111111111111111111111111111111111111111110000"),
("000011000000000111111111100000000000111111111110001111110000"),
("000111000000000001111111100000000000111111110000000001111000"),
("000111000000000000111111100000000000111111100000000000111000"),
("000111000111111000011111100011111111111111000011111110111000"),
("001111000111111100011111100011111111111110000111111111111100"),
("001111000111111100011111100011111111111110001111111111111100"),
("001111000111111100011111100011111111111110001111111111111100"),
("001111000111111100011111100011111111111100011111111111111100"),
("001111000111111000011111100011111111111100011111111111111110"),
("011111000000000000111111100000000001111100011111111111111110"),
("011111000000000011111111100000000001111100011111111111111110"),
("011111000000000011111111100000000001111100011111111111111110"),
("011111000111110001111111100011111111111100011111111111111110"),
("011111000111110000111111100011111111111100011111111111111110"),
("011111000111111000111111100011111111111100001111111111111110"),
("011111000111111000011111100011111111111110001111111111111110"),
("011111000111111100011111100011111111111110000111111111111110"),
("001111000111111100011111100011111111111111000011111110111110"),
("001111000111111110001111100000000000111111100000000000111100"),
("001111000111111110001111100000000000111111110000000001111100"),
("001111000111111111001111100000000000111111111110001111111100"),
("001111111111111111111111111111111111111111111111111111111100"),
("000111111111111111111111111111111111111111111111111111111000"),
("000111111111111111111111111111111111111111111111111111111000"),
("000111111111111111111111111111111111111111111111111111111000"),
("000011111111111111111111111111111111111111111111111111110000"),
("000011111111111111111111111111111111111111111111111111110000"),
("000001111111111111111111111111111111111111111111111111100000"),
("000000111111111111111111111111111111111111111111111111100000"),
("000000111111111111111111111111111111111111111111111111000000"),
("000000011111111111111111111111111111111111111111111110000000"),
("000000001111111111111111111111111111111111111111111100000000"),
("000000000111111111111111111111111111111111111111111000000000"),
("000000000111111111111111111111111111111111111111111000000000"),
("000000000001111111111111111111111111111111111111100000000000"),
("000000000000111111111111111111111111111111111111000000000000"),
("000000000000011111111111111111111111111111111110000000000000"),
("000000000000001111111111111111111111111111111100000000000000"),
("000000000000000011111111111111111111111111110000000000000000"),
("000000000000000000111111111111111111111111000000000000000000"),
("000000000000000000000111111111111111111000000000000000000000"),
("000000000000000000000000011111111110000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000")
);

signal bCoord_X : integer := 0;-- offset from start position 
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';

--		
signal objectEndX : integer;
signal objectEndY : integer;


signal mVGA_R	: std_logic_vector(2 downto 0); --	,	 			//	VGA Red[2:0]
signal mVGA_G	: std_logic_vector(2 downto 0); --	,	 			//	VGA Green[2:0]
signal mVGA_B	:  std_logic_vector(1 downto 0); --	,  				//	VGA Blue[1:0]


begin

-- Calculate object end boundaries
objectEndX	<= object_X_size+StartX;
objectEndY	<= object_Y_size+StartY;

-- Signals drawing_X[Y] are active when obects coordinates are being crossed

-- test if ooCoord is in the rectangle defined by Start and End 
	drawing_X	<= '1' when  ( (oCoord_X  >= StartX) and  (oCoord_X < objectEndX) ) else '0';
    drawing_Y	<= '1' when  ( (oCoord_Y  >= StartY) and  (oCoord_Y < objectEndY) ) else '0';


bCoord_Y <= (oCoord_Y - StartY) when ( (drawing_X = '1') and  drawing_Y = '1'  ) else 0 ; 


process (RESETn, CLK)
  
   begin
	if drawing_Y = '1' then
	bCoord_X <= (oCoord_X - StartX);
		if (drawing_X = '1') then
			bCoord_X <= (oCoord_X - StartX);
		else
			bCoord_X <= 0 ;
		end if;
	end if;
	if RESETn = '0' then
	    mVGA_RGB <=  mVGA_R & mVGA_G &  mVGA_B ;
		-- defining three rectangles 
		mVGA_R <= "000";
		mVGA_G <= "000"; 
		mVGA_B <= "00";
		drawing_request	<=  '0';
		elsif rising_edge(CLK) then
		    mVGA_RGB <=  mVGA_R & mVGA_G &  mVGA_B ;
			-- defining three rectangles
			if(Record1Enable='0') then
				mVGA_R <= "000";
				mVGA_G <= "000"; 
				mVGA_B <= "00";
			else
				mVGA_R <= "111";
				mVGA_G <= "000"; 
				mVGA_B <= "00";
			end if;
			drawing_request	<= drawing_X and drawing_Y and object(bCoord_Y , bCoord_X) ; -- get from mask table if inside rectangle 
	end if;

  end process;

		
end behav;		
		